module assignemt;
integer alpha, beta;

initial begin
    alpha = 4;
    beta = 3;
    beta <= beta + alpha;
    alpha <= alpha + beta;
    alpha = alpha - 1;
    $display("display values Alpha=%0d Beta=%0d", alpha, beta);
end
initial $monitor("Monitor values Alpha=%0d Beta=%0d", alpha,
beta);

endmodule